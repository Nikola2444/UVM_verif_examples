`ifndef TEST_BASE_SV
 `define TEST_BASE_SV

class test_base extends uvm_test;

   calc_env env;
   calc_config cfg;
    
   `uvm_component_utils(test_base)

   function new(string name = "test_base", uvm_component parent = null);
      super.new(name,parent);
   endfunction : new

   function void build_phase(uvm_phase phase);
      super.build_phase(phase);
       cfg = calc_config::type_id::create("cfg");      
       uvm_config_db#(calc_config)::set(this, "env", "calc_config", cfg);      
       env = calc_env::type_id::create("env", this);      
   endfunction : build_phase

   function void end_of_elaboration_phase(uvm_phase phase);
      super.end_of_elaboration_phase(phase);
      uvm_top.print_topology();
   endfunction : end_of_elaboration_phase

    function void init_vseq(virtual_seq vseq);
	vseq.interface1_seqr = env.agent1.seqr;
	vseq.interface2_seqr = env.agent2.seqr;
	vseq.interface3_seqr = env.agent3.seqr;
	vseq.interface4_seqr = env.agent4.seqr;
    endfunction: init_vseq

endclass : test_base

`endif
